CircuitMaker Text
5.6
Probes: 1
Q1_3
Transient Analysis
0 467 426 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 30 100 10
180 79 1274 744
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.412181 0.500000
348 175 1442 449
9961490 0
0
6 Title:
5 Name:
0
0
0
13
9 Resistor~
219 259 255 0 4 5
0 5 2 0 -1
0
0 0 864 90
5 1000k
3 2 38 10
4 HAND
8 -11 36 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
40229.8 3
0
12 SPDT Switch~
164 256 300 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4704 270
0
5 Short
7 -4 42 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
5616 0 0
2
40229.8 2
0
12 SPST Switch~
165 254 342 0 2 11
0 5 4
0
0 0 4704 90
0
5 Touch
1 -6 36 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9323 0 0
2
40229.8 1
0
7 Ground~
168 259 169 0 1 3
0 2
0
0 0 53344 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
317 0 0
2
40229.8 0
0
10 Capacitor~
219 363 476 0 1 5
0 0
0
0 0 832 90
5 100nF
4 0 39 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 16643792
67 0 0 0 1 0 0 0
1 C
3108 0 0
2
40229.8 0
0
2 +V
167 363 142 0 1 3
0 7
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4299 0 0
2
40229.8 0
0
4 LED~
171 465 517 0 2 2
10 13 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9672 0 0
2
40229.8 0
0
13 PNP Darling1~
219 457 391 0 3 7
0 14 3 15
0
0 0 848 692
10 MMBTA63LT1
44 1 114 9
2 Q1
29 -10 43 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 SOT-23
7

0 3 1 2 3 1 2 16594728
88 0 0 256 1 1 0 0
1 Q
7876 0 0
2
40229.8 0
0
7 Ground~
168 465 557 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
5.89466e-315 5.30499e-315
0
7 Ground~
168 363 554 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
5.89466e-315 5.32571e-315
0
2 +V
167 465 152 0 1 3
0 15
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
5.89466e-315 5.38788e-315
0
9 Resistor~
219 363 343 0 4 5
0 4 7 0 1
0
0 0 880 90
5 1000k
6 -1 41 7
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 250
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
40229.8 0
0
9 Resistor~
219 465 463 0 2 5
0 13 14
0
0 0 880 90
3 100
6 0 27 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7678 0 0
2
40229.8 0
0
13
0 3 2 0 0 0 0 0 2 3 0 3
259 227
251 227
251 284
2 0 4 0 0 16 0 3 0 0 7 3
255 358
255 391
363 391
1 2 2 0 0 0 0 4 1 0 0 2
259 177
259 237
1 1 5 0 0 0 0 2 3 0 0 2
255 318
255 324
1 2 5 0 0 0 6 1 2 0 0 4
259 273
259 286
259 286
259 284
1 2 7 0 0 12416 0 6 12 0 0 2
363 151
363 325
1 0 4 0 0 0 0 12 0 0 10 2
363 361
363 391
2 1 2 0 0 128 0 7 9 0 0 2
465 527
465 551
1 1 13 0 0 4224 0 13 7 0 0 2
465 481
465 507
2 2 4 0 0 4224 0 5 8 0 0 3
363 467
363 391
433 391
1 2 14 0 0 20608 0 8 13 0 0 2
465 413
465 445
1 3 15 0 0 28800 0 11 8 0 0 2
465 161
465 369
1 1 2 0 0 12416 0 10 5 0 0 2
363 548
363 485
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
