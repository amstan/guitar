CircuitMaker Text
5.6
Probes: 1
Q1_1
Transient Analysis
0 466 287 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
180 79 1274 744
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.412181 0.500000
348 175 1442 449
9961490 0
0
6 Title:
5 Name:
0
0
0
15
2 +V
167 417 140 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5130 0 0
2
40229.8 0
0
4 LED~
171 465 200 0 2 2
10 8 5
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
391 0 0
2
5.89466e-315 0
0
10 Capacitor~
219 363 413 0 2 5
0 2 7
0
0 0 848 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 250
67 0 0 0 1 0 0 0
1 C
3124 0 0
2
5.89466e-315 0
0
12 NPN Trans:B~
219 411 367 0 3 7
0 4 7 9
0
0 0 848 0
3 NPN
17 0 38 8
2 Q2
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3421 0 0
2
5.89466e-315 5.26354e-315
0
7 Ground~
168 465 457 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
5.89466e-315 5.30499e-315
0
7 Ground~
168 363 451 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
5.89466e-315 5.32571e-315
0
12 SPST Switch~
165 362 286 0 10 11
0 12 12 0 0 0 0 0 0 0
1
0
0 0 4720 90
0
2 S2
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8901 0 0
2
5.89466e-315 5.34643e-315
0
2 +V
167 367 153 0 1 3
0 10
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89466e-315 5.3568e-315
0
12 SPDT Switch~
164 364 244 0 10 11
0 12 12 10 0 0 0 0 0 0
1
0
0 0 4720 270
0
2 S1
9 -4 23 4
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4747 0 0
2
5.89466e-315 5.36716e-315
0
12 NPN Trans:B~
219 460 391 0 3 7
0 6 9 2
0
0 0 848 0
3 NPN
17 0 38 8
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
972 0 0
2
5.89466e-315 5.37752e-315
0
2 +V
167 465 152 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.89466e-315 5.38788e-315
0
9 Resistor~
219 416 238 0 4 5
0 4 3 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 16600452
82 0 0 0 1 0 0 0
1 R
9998 0 0
2
40229.8 0
0
9 Resistor~
219 465 250 0 2 5
0 6 5
0
0 0 880 90
3 100
6 0 27 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3536 0 0
2
40229.8 0
0
9 Resistor~
219 363 326 0 2 5
0 7 12
0
0 0 880 90
4 100k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 16718392
82 0 0 0 1 0 0 0
1 R
4597 0 0
2
5.89466e-315 5.39306e-315
0
9 Resistor~
219 367 199 0 4 5
0 12 10 0 1
0
0 0 880 90
5 1000k
-2 0 33 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 16595128
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
5.89466e-315 5.39824e-315
0
15
1 2 3 0 0 4224 0 1 12 0 0 4
417 149
417 219
416 219
416 220
1 1 4 0 0 4224 0 12 4 0 0 2
416 256
416 349
2 2 5 0 0 4224 0 2 13 0 0 2
465 210
465 232
1 1 6 0 0 4224 0 13 10 0 0 2
465 268
465 373
3 1 2 0 0 4224 0 10 5 0 0 2
465 409
465 451
0 2 7 0 0 4096 0 0 4 10 0 4
363 367
403 367
403 367
393 367
1 1 8 0 0 4224 0 11 2 0 0 2
465 161
465 190
3 2 9 0 0 8320 0 4 10 0 0 3
416 385
416 391
442 391
0 3 10 0 0 8320 0 0 9 13 0 3
367 171
359 171
359 228
1 2 7 0 0 4224 0 14 3 0 0 2
363 344
363 404
2 2 12 0 0 4224 11 7 14 0 0 2
363 302
363 308
1 1 2 0 0 0 0 6 3 0 0 2
363 445
363 422
1 2 10 0 0 0 0 8 15 0 0 2
367 162
367 181
1 1 12 0 0 4224 0 9 7 0 0 2
363 262
363 268
1 2 12 0 0 4224 13 15 9 0 0 4
367 217
367 230
367 230
367 228
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
