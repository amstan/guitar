CircuitMaker Text
5.6
Probes: 1
r1[i]
Operating Point
0 672 374 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
340 170 30 100 10
344 81 1278 648
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
512 177 1446 460
9961490 0
0
6 Title:
5 Name:
0
0
0
12
2 +V
167 884 299 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9172 0 0
2
40232 2
0
7 Ground~
168 884 514 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7100 0 0
2
40232 1
0
4 LED~
171 884 456 0 2 2
13 3 2
0
0 0 880 0
4 LED3
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3820 0 0
2
40232 0
0
2 +V
167 781 302 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7678 0 0
2
40232 2
0
7 Ground~
168 781 517 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
961 0 0
2
40232 1
0
4 LED~
171 781 459 0 2 2
12 5 2
0
0 0 880 0
4 LED2
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3178 0 0
2
40232 0
0
4 LED~
171 673 461 0 2 2
10 7 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3409 0 0
2
40232 0
0
7 Ground~
168 673 519 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3951 0 0
2
40232 0
0
2 +V
167 673 304 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8885 0 0
2
40232 0
0
9 Resistor~
219 884 384 0 4 5
0 3 4 0 1
0
0 0 880 90
2 82
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
40232 3
0
9 Resistor~
219 781 387 0 4 5
0 5 6 0 1
0
0 0 880 90
3 150
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
40232 3
0
9 Resistor~
219 673 389 0 4 5
0 7 8 0 1
0
0 0 880 90
3 180
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 16687748
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
40232 0
0
9
2 1 2 0 0 4240 0 3 2 0 0 2
884 466
884 508
1 1 3 0 0 4240 0 10 3 0 0 2
884 402
884 446
2 1 4 0 0 4240 0 10 1 0 0 2
884 366
884 308
2 1 2 0 0 0 0 6 5 0 0 2
781 469
781 511
1 1 5 0 0 4224 0 11 6 0 0 2
781 405
781 449
2 1 6 0 0 4224 0 11 4 0 0 2
781 369
781 311
2 1 2 0 0 128 0 7 8 0 0 2
673 471
673 513
1 1 7 0 0 4224 0 12 7 0 0 2
673 407
673 451
2 1 8 0 0 4224 0 12 9 0 0 2
673 371
673 313
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
